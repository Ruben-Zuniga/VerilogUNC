module count (

    output              valid,
    input       [2:0]   i_sw,
    input               i_reset,
    input               clock

);



endmodule