module led_project(

    input       [3:0]   i_sw,
    input               i_reset,
    input               clock,
    output      [3:0]   o_led,
    output      [3:0]   o_led_b,
    output      [3:0]   o_led_g
    
);

endmodule